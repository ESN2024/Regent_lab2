
module lab2_sys (
	clk_clk,
	pio_0_seg_export,
	reset_reset_n);	

	input		clk_clk;
	output	[11:0]	pio_0_seg_export;
	input		reset_reset_n;
endmodule
